module xorr (input din1, din2, output dout);

assign dout = din1 ^ din2;

endmodule
